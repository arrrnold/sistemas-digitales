----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:58:49 11/23/2021 
-- Design Name: 
-- Module Name:    MUX4bitsPROCESS - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

				entity CONC4bits is
					 Port ( A0 : in  STD_LOGIC;
							  A1 : in  STD_LOGIC;
							  A2 : in  STD_LOGIC;
							  A3 : in  STD_LOGIC;
							  control : in  STD_LOGIC_VECTOR (1 downto 0);
							  salida : out  STD_LOGIC);
				end CONC4bits;

				architecture Behavioral of CONC4bits is
				begin

					 process (A0,A1,A2,A3,control)
					 begin

						  salida <=   A0 when (control="00") else
										  A1 when (control="01") else
										  A2 when (control="10") else
										  A3 when (control="11") else
										  0;
					 end process;


				end Behavioral;



